`timescale 1ns / 1 ps

// 16 x oversample

module baud_rate_generator #(parameter oversample=0)
(
   input         clk_i,
   input         rst_i,
   output        rx_tick_o,
   output        tx_tick_o,
   input  [15:0] baud_div_i 
);
    
   reg rx_tick_o_r ;
   reg tx_tick_o_r ;
   
   assign rx_tick_o = rx_tick_o_r;
   assign tx_tick_o = tx_tick_o_r;
       
   wire [15:0] max_r_clock;
   wire [15:0] max_t_clock;
   assign max_r_clock = baud_div_i >> (oversample == 5'd16 ? 3'd4 : oversample == 4'd8 ? 2'd3 : 0);
   assign max_t_clock = baud_div_i;
   
   reg [15:0] rx_counter ;
   reg [15:0] tx_counter ;

   always @(posedge clk_i) begin
 
      if(!rst_i) begin // rst_i == 0 ise resetlenecek
         rx_counter  <= 32'd0;
         rx_tick_o_r <= 1'b0;
         tx_counter  <= 32'd0;
         tx_tick_o_r <= 1'b0;
      end
      
      else begin 
      
         // rx clock
         
         if (rx_counter == (max_r_clock-1'b1)) begin
            rx_counter  <= 32'd0;
            rx_tick_o_r <= 1'b1;
         end 
         else if (rx_counter > (max_r_clock-1'b1)) begin
            rx_counter  <= 32'd0;
            rx_tick_o_r <= 1'b0;
         end
         else begin
            rx_counter  <= rx_counter + 1'b1;
            rx_tick_o_r <= 1'b0;
         end
         
         // tx clock
         
         if (tx_counter == (max_t_clock-1'b1)) begin
            tx_counter  <= 32'd0;
            tx_tick_o_r <= 1'b1;
         end 
         else if (tx_counter > (max_t_clock-1'b1)) begin
            tx_counter  <= 32'd0;
            tx_tick_o_r <= 1'b0;
         end
         else begin
            tx_counter  <= tx_counter + 1'b1;
            tx_tick_o_r <= 1'b0;
         end
      end
    end
    
endmodule
